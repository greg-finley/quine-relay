module QR;initial begin $write("%s",("let s=(\"Module QR:Sub Main():Dim c,n,s As Object=System.Console.OpenStandardOutput(),t()As Short={26,34,85,127,144,153,196}:For Each c in\\\"BasmCBBBCRE`F<<<<C<`C<B`BBD#CXwasi_snapshot_preview1Jfd_writeBBEEDCDGECB@IUDHmemoryDBH_startBDL|DRBAC BAJlACA4RB9MiCD<AERCA>D!BE@ABRCABRCABRCAJ!CE@ B-BB CACk:CvACqRC COBMADRCACRCADRCABRCABRC BACj:B-BBOBMADRCADRCADRCAFRCMM}CBABM~(BBBCBBB,BBBDBBB0BBBDBBB4BBB=BBB?BBB;BBB ...\\\\t..\\\\n..(module(import:wasi_snapshot_preview1::fd_write:(func(param i32 i32 i32 i32)(result i32)))(memory(export:memory:)(data :\\\\08\\\\00\\\\00\\\\00$:))(func(export:_start:)i32.const 1 i32.const 0 i32.const 1 i32.const 0 call 0 drop))\\\":c=Asc(c):If c=36:For c=0To 11:s.WriteByte(If(c Mod 3,Asc(607043.ToString(\\\"x8\\\")(1Xor 7-c*2\\\\3)),92)):Next:Else:n=(c>12"));
$write("%s",("4)*(8*c-39229):Do While n>127:s.WriteByte(128+(127And n)):n\\\\=128:Loop:s.WriteByte(If(c<125,If((c-1)\\\\7-8,c+66*(c>65And c<91),t(c-57)),n)):End If:Next:For Each c in\\\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[sub f(s$,n)print(s$);:for i=1to n print(\\\"\\\"\\\\\\\\\\\"\\\");:next:end sub:f(\\\"\\\"write,format=\\\\\\\"\\\"%s%s%s%s\\\\\\\"\\\",\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"write{-}{txt}{echo -E $'(\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put(\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans B(Buffer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans O(n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Chara"));
$write("%s",("cter\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"B:add(Byte(+ 128 n))\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans f(v n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(+(/ n 64)107)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(n:mod 64)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O v\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans D(n)\\\"\\\",2):f(\\\"\\\"{if(< n 4)\\\"\\\",2):f(\\\"\\\"{f(+(* 6 n)9)48\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{if(n:odd-p)\\\"\\\",2):f(\\\"\\\"{D(- n 3)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 27 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f("));
$write("%s",("\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 36 11\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{D(/ n 2)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 21 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 48 20\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans S(Buffer\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"2\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR160,c:=b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR165,t:=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class QR\\\"\\\",2):f(\\\"\\\"{public static void main(String[]a)\\\"\\\",2):f(\\\"\\\"{a=("));
$write("%s",("\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"write(\\\"\\\",4):f(\\\"\\\"'implement main0()=print(^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"BEGIN\\\"\\\",2):f(\\\"\\\"{print(^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"echo ^1^\\\"\\\",4):f(\\\"\\\"'f(s)\\\"\\\",2):f(\\\"\\\"{System.out.print(s);\\\"\\\",2):f(\\\"\\\"}s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"389**6+44*6+00p45*,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(c:(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<stdio.h>^8^nchar*p=(^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Ra#include<iostream>^16^nint main()\\\"\\\",2):f(\\\"\\\"{std::cout<<(^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class Program\\\"\\\",2):f(\\\"\\\"{public static void M83abbSystem.Console.Write(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Quine Relay Coffee.^64^n^64^nIngredients.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=9;i++<126;)[3pva$^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"} g caffeine \\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}I3b54rja^64^nMethodv4f#aeach(char c in(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\"));
$write("%s",("\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")))^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2al3dp3c[2cs3c,3l[2k@3kqa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")s rts(ecalper.h3eja^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"     53c4a SUTATS(egassem^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"rts(nltnirp(])]^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NUR POTSu4cba.C3dh3dX3bba[65bX4df5lga\\\"\\\",2):f(\\\"\\\"};)06xm3f$3loa)1(f\\\"\\\",2):f(\\\"\\\"{#qp]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\"));
$write("%s",("\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[p]#3sv3r23)ga3(f\\\"\\\",2):f(\\\"\\\"{#.33)ba7g4-ba5R4w23F&7d33&q7u53sda,4353.ma^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' D ; EYB RCL4/v4+ja13(f\\\"\\\",2):f(\\\"\\\"{#DNEm4[m4ada. A~5[p"));
$write("%s",("4deaPOTSn4[#5e~5[o4boaRQ margorp dnex4[x4abaS*5[m4c2<[ba9i4[i4dba&#6[k4agaS POOL&<[77dba^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'j4[j4[j4gda&,)(6[<>cga. TNUO<7[s4bfa(rahcf:[(5dgaB OD 0?>[t4cca&,+<[ha9(f\\\"\\\",2):f(\\\"\\\"{#)A26[9=d4=[,6cqaEUNITNOC      01z4[a9c,5[U8dJ7[WFeeaRC .p4[p4aka,1=I 01 ODt4[OKecaPUq4[*I[5<gva;TIUQ;)s(maertSesolC;dYe$4Rra322(f\\\"\\\",2):f(\\\"\\\"{#tiuqn\\\"\\\",2):f(\\\"\\\"})652=5[qa^32^\\\"\\\",2):f(\\\"\\\"})974(f\\\"\\\",2):f(\\\"\\\"{#n\\\"\\\",2):f(\\\"\\\"})215iY3b8,ya99(f\\\"\\\",2):f(\\\"\\\"{#etalpmetdne.n\\\"\\\",2):f(\\\"\\\"})4208[.zX3ca02-Y[v3bda116~K[-L[j4ldamif+6[ga)30341\\\"\\\",2):f(\\\"\\\"}5[,6[j4l"));
$write("%s",("bat(6[(6c%a315133A71/129@31916G21661421553/04[04c(a%%%%\\\"\\\",2):f(\\\"\\\"}*+1%%%%811 -\\\"\\\",2):f(\\\"\\\"})48361(f\\\"\\\",2):f(\\\"\\\"{#j:+1 j@34[34cbawm4[m4cl4[l4cbaWm4[m4cba\\\"\\\",2):f(\\\"\\\"{m4[m4cva)(esolc.z;)][etyb sa)t=[#>[j4[~Jjca69m4[x5[j4lba,l4[w5[j4hla!\\\"\\\",2):f(\\\"\\\"})23(f\\\"\\\",2):f(\\\"\\\"{#~~v4[%5[j4hea(rt.o4[z5[j4hba)A7dda\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};l3efa~~dneo3hra~~~~PUEVIGESAELPnr3ala~~1,TUODAERw3a63j$a(etirw;\\\"\\\",2):f(\\\"\\\"};u=:c;))652%%%%)u-c((||13jda#-<q3jda||i)3mhaBUS1,ODs4qka)3/4%%%%i(N4cx5kU4xPa2=:/t;2%%%%t+2*u=:u\\\"\\\",2):f(\\\"\\\"{od7 ot0 yreve;i-=:u;1=:+i\\\"\\\",2):f(\\\"\\\"{od))1(evom(dro=:t elihw?s;)s*45oi5vv3jd7dladohtem dne.s3dganrutern3d~aV);gnirtS/gnal/avajL(nltnirp/+Za|atnirP/oi/avaj lautrivekovniJ3d.4j[2cib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\"\\\",2):f(\\\"\\\"{)0>2%%%%++i(fi;48%%%%)31-)i>3c&as(+87*q=q\\\"\\\",2):f(\\\"\\\"{);68312<i;(rof;n)rahc(+K4r[2k*3&oa=]n[c);621<n++r4aqa0=q,0=n,0=i tni;N3&bc6ayi4asdRbQehlxfvfalRf<bedRb;fkW;agb-a|dzdxdRfGb8aqeRdYd5a4<Gi;agb-epb>aqeRdHa>aJaRaAdteFbaeIfOa5aac2gb26f9azb<a4aLa7a;a4a<aPhhmkdxd;aNa?c6a|eebHaFaIaebzeJaeb9a/a6a2dQbUe-f2a-I3bga5d6cRbE3gYc-f/aof0fRfkh9kEf.b2e6aRa;d6sogB\\\"\\\",2):f(\\\"\\\"{Gh;aTapc4aLcEeyiof6amc<byg-f?lsbvhgUWfybxcxcAUUeAa2a6a\\\"\\\",2):f(\\\"\\\"}g7a6a@a\\\"\\\",2):f(\\\"\\\"{g:a?aMbKaKa6a?e:a@aEa2a|gZfMbbgli>a:b1a-gfmUf\\\"\\\",2):f(\\\"\\\"{bHa4atc3b3+rI0qrIEcZFJaMa\\\"\\\",2):f(\\\"\\\"}bJaZzEc-bJaJaUa-bJaMdJa8bq2;a+wTaKa+wTaQA1j\\\"\\\",2):f(\\\"\\\"}bKRSaSaNa+b9bKa+wA|Ta+w+wTa8bNa+bm\\\"\\\",2):f(\\\"\\\"}JaLaJa8bN;N"));
$write("%s",("an4c\\\"\\\",2):f(\\\"\\\"{3ava3++b:b0qrI0q+b1j\\\"\\\",2):f(\\\"\\\"}bJaH/3a=3b-aHaJaFdo5;a+wUa:aUa:aq2viSfQfGl4airsbsb2be3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'maviDa-a|bf>-aF6asacKUe>a5j\\\"\\\",2):f(\\\"\\\"{gKaKa|gZf(6cgaagQjkg,6esasbvh*b-a/bxcHa|fDke3c4c\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"{gph\\\"\\\",2):f(\\\"\\\"{gvg1a-g\\\"\\\",2):f(\\\"\\\"{bHaDkRf-e:a:a\\\"\\\",2):f(\\\"\\\"}bHa?a\\\"\\\",2):f(\\\"\\\"{gJa\\\"\\\",2):f(\\\"\\\"}b5aAdte@a1a-g0iDkxcpb7anb2b:b\\\"\\\",2):f(\\\"\\\"{g2f@j@d-aIfekxcHa>a1a-gigggti-aUf0ixiRf-f-gSf|fDkzeSgxiHack;a/aDh<b+hWh<apb/aDhWhnblK7b:b\\\"\\\",2):f(\\\"\\\"{g/aDh-f-g+gFa,i|b1ali3b:b\\\"\\\",2):f(\\\"\\\"{g9hHaDkHaUe-iCe|bx"));
$write("%s",("c3b0a:b\\\"\\\",2):f(\\\"\\\"{gIa|bzeJa|g5buaQbxi<b=a-a=m*c3bxdUem3aea|b9ai3eta2bMa7arh|bphnhlhjh9m3hAaAd\\\"\\\",2):f(\\\"\\\"}4PcgfvfOhJh7aEa|b0k.kMa=m*cEc,dJa>a2aIfzjMgMa=m|b<i+cbi6a13iYa|b<iV?2t8g/aDh=apiRaWJCdlbaq6,Hwpiak6a7b5ackRfwb\\\"\\\",2):f(\\\"\\\"}jUe2b5a9gYigFhcfsOiOiOu0c/bxd;a<hoj3?aea6a2bZ>ekc8DCL6a\\\"\\\",2):f(\\\"\\\"}n2a5ajn@J\\\"\\\",2):f(\\\"\\\"}g6hjkavOi6aUhinHa1dmdLhRfWkLkHa:eWkLk0l<b3bxd6aIh8kPh\\\"\\\",2):f(\\\"\\\"}l/SkivftfTF;aXiccoJpbD6tvZbrpnbpgujsjiih0RiVkuhTk4j<b<b<bFj:b<j<b<b,cKjHj.MKjEa;k*k,cCjMi9a+Y-agJ,b,cKj=a9a7bubxbs3e13ecaCj13gA3a13kgaJb7bdgo3eka;p?au.9av2)3cmakirkpj7k,cKji3asa-aJd8Cfh,cKjsbHa\\\"\\\",2):f(\\\"\\\"}gw5ciaVjDjCaLi46aka7jhk4j<bzeCCc/3gda2k3m3fKa<kLi6a<bkicjQ\\\"\\\",2):f(\\\"\\\"}0>8R>L2a2a=HekOk0iwb\\\"\\\",2):f(\\\"\\\"}jRf@a>anc:e7b5aWf=anbekybvk5a,bJa6acAa%aub9h5aUgwb"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"}jHa:e-b9a9b9a2kekyg>am3a\\\"\\\",2):f(\\\"\\\"{a@a@aekyg@a>a:a|b9a0b9a@a>aLBakb>e|bPg9bJa0bekyg-b9a2k9aCaAaJa9beknbJa6a|b5a,bRf:e-b0kwN-ajh9apb2lDL6Vvi=Hyg8bAdGh-a=H+3bb-a=Hyg7s3h13albXb;d9f/bxd6a-b9a8b9a7bJcJayb>a;pki>aJa*c@dxc?b,b0G>aJa-b>lteUe@a;M2b5aDci>:atcJaub5aEcxbh0,bgFJaUgu7eeaJkHkq;e^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'cSkQkpb;awb\\\"\\\",2):f(\\\"\\\"}jslx\\\"\\\",2):f(\\\"\\\"{0>8R7V@TuZ4@sZJdHdSl1nqn8lbm-n+nwnR>0nhc/*5C|xu+<4pxnx\\\"\\\",2):f(\\\"\\\"{|MwPEMwfr|x=Xl/FAt4lb.bcJV4Cap+zvl5UG2u.b6\\\"\\\",2):f(\\\"\\\"}aoroirM4fr1\\\"\\\",2):f(\\\"\\\"{-bGnss6b1bgb+oZas0U8kYt>DoSat03G2bgbO0qp.qu"));
$write("%s",("u?aG/Q86b1b\\\"\\\",2):f(\\\"\\\"}pE7Ea/8.yhb.u/Kt4hbso2h0b.<k5cydvb+:Tp?o>-bb?9q-+dhr96bywtCatQVmt46Jeb9\\\"\\\",2):f(\\\"\\\"{XQB>cR?\\\"\\\",2):f(\\\"\\\"}yw|ba0wopLhjT\\\"\\\",2):f(\\\"\\\"{WOTpo\\\"\\\",2):f(\\\"\\\"}u/4Xab.00-q*Damu61-s4J1xgJYavb;qlb8o\\\"\\\",2):f(\\\"\\\"{59H23Dq+w9-zb\\\"\\\",2):f(\\\"\\\"{bTpYnVC+ww+-=Kp6AyF2bWaBaJZBaZpkiBlio.02|f7CacbpD=\\\"\\\",2):f(\\\"\\\"{cba5FVV|ybZnP;\\\"\\\",2):f(\\\"\\\"{b.q?\\\"\\\",2):f(\\\"\\\"},C7b|TWncKDQEa+FyJ/*-bav>rK2Y,8/mb-bibt4-Jz0.b0LXn*bkr-J@oYimQ|*K-OAMq7bV7hwXQ3:u6Ww\\\"\\\",2):f(\\\"\\\"}K\\\"\\\",2):f(\\\"\\\"{OP|\\\"\\\",2):f(\\\"\\\"{b5py&6f&d4b,bCq\\\"\\\",2):f(\\\"\\\"}sXakbRBMKjbm|<aZhebEaCay0a0u;A9jwSau:wtWaVaFSFr2L\\\"\\\",2):f(\\\"\\\"}59zCrH=Q>nyWp/r00a\\\"\\\",2):f(\\\"\\\"{Kv*VV*/6+9>aIu|wLW=ogbNtZaibY\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{6o/nX<I7qa/Ui1;sqivEaYrUn5bDargF4BaEa5b7urL:oBaOwg@XKAa+tZaxSP2AaYav3tby"));
$write("%s",("9Hx2|*;a6h@mHe\\\"\\\",2):f(\\\"\\\"{/|/yC9lbSakiTTBaEaiogoUAooPaMRPq>a3H:Tdbhb6bX|96BaEa-bAaZ0-s@RF|nox@jo0odPg@2Fetu6oo-;W,3|>a4b,bTAPa.6e%czbSPzbz@d,SaVvoT/bLR3bP8\\\"\\\",2):f(\\\"\\\"{6qRoRooTaI-Ta3|y6lIfReSa*cR9rTaEa3:@qPPyPqFYWjb-2DarxM|9b=aYWjbo?hAVaFA5-0-uj,v,v4|PP1-6p6F,b@a0-m6qqB|4|By,bl5-2ONKxaQh@v0U\\\"\\\",2):f(\\\"\\\"{5G|Qlbhbb7N;-bbo0rl5CEQa9rMw3:-p+2P96p,\\\"\\\",2):f(\\\"\\\"{L;+bl5.b,bbohb9tO3aVa.bj9fTSam+9r59-Shy3:Ta.b3qws8yEaBabXDa,bbDgbrxCas7z2gbjb*rboUGDad\\\"\\\",2):f(\\\"\\\"}CvlbUGDaHrCx9A1Y9fFbgbHrub7|eb3,-Pz9=2ubDa31*by9K>tbqq1V//@qhbPp-bSt=\\\"\\\",2):f(\\\"\\\"{kP<on-h\\\"\\\",2):f(\\\"\\\"}hb*rz@?ey0p<DT/*7b6+dbhb;<WOWaOp0b+o\\\"\\\",2):f(\\\"\\\"}o:o2blCTaE2vbC?\\\"\\\",2):f(\\\"\\\"{OC?J|tbRp<kDa\\\"\\\",2):f(\\\"\\\"{OC?lCLp\\\"\\\",2):f(\\\"\\\"{K=shbq<DaiFu*3:/*hb#3c4bZ5t06b8oJLWaaxhblb-bOahbvre1q<Dap|<aD"));
$write("%s",("aabzO-wTaiVWAib7bEaUpVruB.FvbYxF0cO@1q8Yha6ON?9LNJN|bHNffEN2TL54b/QD5d|9ouSBakGCaBnh*mbUa,hUoxbeN[9gOaTao>Pa=a5o8N.*\\\"\\\",2):f(\\\"\\\"{btbOjibBaRahbhbq3.GS<F5Ravb+o.*f0az=ayxSB1b<sHpH.q<17<aVv-bi3a4byPBP6oc\\\"\\\",2):f(\\\"\\\"}34/ux:n-0.hbAqkiLVlbCa79W-DaYt>7?.6oOaPa1Mmu=8vQ*6buEOub=a84/bYwy\\\"\\\",2):f(\\\"\\\"}t<w,?a9bDauyQaFwAa9bc|=,iCBaB4UXzbN,K38wC0sIgb3*40;7lz,tC5L,S3Wka<N:BDL6VddY3kfduEKh1A>-tbVa3Hkb4.q*k5Eu*|Wa:rxbcKuSx*FJlb37S,bb|Hcbvpkr2bcoa\\\"\\\",2):f(\\\"\\\"{0|tbHrybiOS,qr/uo3S2qqPsaBCq6F\\\"\\\",2):f(\\\"\\\"}.tb=wHpk=psuBzb>U7<lqt@tbv9mFNx8gIhVa+b.d=sX+4ATAtbFayxl\\\"\\\",2):f(\\\"\\\"{uP5.AaX3Yaf2AaJ8kyWi@z3yWi6--brR3T1T-b2t<>mYTMccUoxbv+1bTAtbWD4bDp\\\"\\\",2):f(\\\"\\\"{+IZVw@*TaV;zPbb-ZZtbFI|ir@*Oyhvw>3ba6qy*bX1<\\\"\\\",2):f(\\\"\\\"}YN-iU9eKafrutjbpUbcibfbwT.E?azbY,hP:T1|yTabPPNadPjb\\\"\\\","));
$write("%s",("2):f(\\\"\\\"}LpsebV6W*RPH+O\\\"\\\",2):f(\\\"\\\"{89D3X7XR1Ajbj4a/cj3tb-F8o\\\"\\\",2):f(\\\"\\\"{4RalwGH4bd4qit8Ss|@<kkiErCrAr?rYNd,L\\\"\\\",2):f(\\\"\\\"{+9ib0LrRhjmb6bhA?airx,Xi/|\\\"\\\",2):f(\\\"\\\"{bMS|bpOU*jBwbXC\\\"\\\",2):f(\\\"\\\"}Gf<L|01S?7bebU83zcOO18o-zvuItyF5wK->az4|btjFgsqIwhbg,L2BF17MmzbRFmbEGWr:T:-hbJ88oQvbb5E6zPaybWiZ|pD,b,HUi*6kb;TDnQa5\\\"\\\",2):f(\\\"\\\"}+V96Ca;>wv,6ecacbl4bkd|Y,FU:s:-/rkrzqEafbfbcReb9y:-hbXXG/eb1bn\\\"\\\",2):f(\\\"\\\"{:fgJ@.jQA3z/l67b8oNaw,u,hZ8**;5,>qPaSG>*xLu*zTl/*3kbF|XpH+;<rXOIbEebiOSaZaJx*u6q+b2b@QGspp\\\"\\\",2):f(\\\"\\\"}b/|?|MV*+q*>v=t|*bqJhG-ExKSd/y8/OvXX11\\\"\\\",2):f(\\\"\\\"{ib1;8bY/tY1tz\\\"\\\",2):f(\\\"\\\"}c;Xs?0BaNCu@p3XM01b*0ul6Sawb|@Val/0bViO1:\\\"\\\",2):f(\\\"\\\"{O7B*\\\"\\\",2):f(\\\"\\\"}b<s.xPsabcqb7j>Q@iRqq*uyxcBtr-bavWa0B=Hk=a6bBbQJB/Y/HI@,<@yPvXO1zbss95ITgvHz+v8bdbZasJEw;*1\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"{x6Ty=XcMzb:Q.+lzazyuzrlzaz7b64Pa\\\"\\\",2):f(\\\"\\\"{tr*i=:\\\"\\\",2):f(\\\"\\\"{R>cyNLPa\\\"\\\",2):f(\\\"\\\"}*n+sp=aUaJvSytbvAd4ezWqorNau;hw-K:,3b8,A3a0byuV\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"plzaz\\\"\\\",2):f(\\\"\\\"{typ/ytbV+UaaQYIlQ\\\"\\\",2):f(\\\"\\\"{9>Olz?G,62Q@,QMB|KS4Bbqfbm@\\\"\\\",2):f(\\\"\\\"}G<1u:RJx8Fr>O7vQ1O1j3XXAXw>8<cbQa,\\\"\\\",2):f(\\\"\\\"}a\\\"\\\",2):f(\\\"\\\"{X5Ba\\\"\\\",2):f(\\\"\\\"}byJAykrUs|RcyNLB\\\"\\\",2):f(\\\"\\\"{kymIXXG/|r3qDybEr6c~d\\\"\\\",2):f(\\\"\\\"}Xz9okyxcB\\\"\\\",2):f(\\\"\\\"{bki*pfb4*.pEp0\\\"\\\",2):f(\\\"\\\"{FAN6ItvbzP@sky>Oeq;qai>azbWaSs/ww>vp;*F+3bPQ?vQ0bqK|UIPp@|6L3P\\\"\\\",2):f(\\\"\\\"}j*3l;mbxr|@\\\"\\\",2):f(\\\"\\\"}*0MTXeVDxwbBqYa@qM0FgibSw@@6,Wa7bc46bzrbyS4tb*be>mbDa;4ebwOPou*i;RFdyss<>,8Va9zD3Zn?amI+b24SGV3Fy6F7b.raxNrybkiy-fR5N\\\"\\\",2):f(\\\"\\\"{bRaz6VCC0zb8o-bmbDqq73hC:fr5.NqDa3Z?|q<-qg1<EpO<Eio|bfbSa|bXaf1vr"));
$write("%s",("+dbYu>PJfxdq*.Q8FqVJCw,vWa0?S=0b0b;+=wa>Y5MseVbbn6MFkt0beTYax\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{Ovptbl9Fn/*Px8uHzBpUatb-99+kbPQNaXwy3VCJQr7tby4u6bbB?6bX\\\"\\\",2):f(\\\"\\\"{4b2QYlVJa6tpHgXrl\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{bH5F5EaLnlbxI8:go4bXrbEuQbEx|?uVJ*Vi>S-WaL;@,6F@a7bh,Q/fox.\\\"\\\",2):f(\\\"\\\"{tjb1<UwD-l/LI?|Va@|hw,Q>-Pa@abrUa2bQHTBkHaOTwl\\\"\\\",2):f(\\\"\\\"{6LYt86PaLh?|VaiJpoEOubXakH753h>xWaPambezhbvsj4Ea@FJfwcK;m?XQH>bbTaO\\\"\\\",2):f(\\\"\\\"{SambyxU8FajBiqWaasIpGaDQBfGafTRBQcR;gbTabbSabbazIzf=BUt@CrEagbQ3|b3J,b-bp<5G*zkb.GiqWaZadbnuUq8y|z\\\"\\\",2):f(\\\"\\\"}vnpav8v9Tnp\\\"\\\",2):f(\\\"\\\"{b<98:go|b@aBaQa8\\\"\\\",2):f(\\\"\\\"{uR-0.1jBw@abJR?hHF|bv552Ao\\\"\\\",2):f(\\\"\\\"{KRBmvITCsw@dwPF@i/bGahSyb1t?9cgbIoJZXwVaG58oC0YazNi>w0p4Xa\\\"\\\",2):f(\\\"\\\"}AnGExS|mbg1tWiy79I8H|VsKu30@U4<FxB9Zslb/b8o-b?H3IX4lEmO"));
$write("%s",("uu17qNq69bD26fPbhof|e\\\"\\\",2):f(\\\"\\\"}1z1zzb\\\"\\\",2):f(\\\"\\\"}IUw\\\"\\\",2):f(\\\"\\\"}IUwAz.pkbq*7vUwdoaQ\\\"\\\",2):f(\\\"\\\"{brg\\\"\\\",2):f(\\\"\\\"{EhCiv,\\\"\\\",2):f(\\\"\\\"{Ba\\\"\\\",2):f(\\\"\\\"}b-bX5tQ\\\"\\\",2):f(\\\"\\\"}*N,Qaf>3v7btQvuCpwBy0Wa=qVaq/LI\\\"\\\",2):f(\\\"\\\"{ysBq7Aaw@mI9Hu6etJQ0z7.MO45CaVaO.YaUA:-Oa=*nxNaEazW4bd/RoevGa.S|3Fajdi,+3a8bLvO|Oa0z\\\"\\\",2):f(\\\"\\\"}bhb?a8/pL@ZwbYaRAE/E0cbSaZrbqgtyvQa/-Ga.SVakbG26vUwVn>yb|Oatba0Oa|baqCSR>NaEaNrPal=L;BnWaRaibREzbmbSayw2b0YAa1tNaabk-Qaj4s<NC868o:6edb@aB,3+89vX4VcoXwTCf\\\"\\\",2):f(\\\"\\\"{S@4SvXs6mb+ICwi>?N*y,rD0K32b\\\"\\\",2):f(\\\"\\\"}8\\\"\\\",2):f(\\\"\\\"}b<1|w0Y0|jx*Ekvj@Ua8t.bGv|*<a:u\\\"\\\",2):f(\\\"\\\"{buRr@>r#3c.bdbyxA-49ZQ,wdbd,|xu-ubFaXalWrITaOTAqqNvqKOM?xt+b\\\"\\\",2):f(\\\"\\\"}bcbM?tAiRWadbvsubFaps@ggJbQfT\\\"\\\",2):f(\\\"\\\"{bB*TqUa?Nh*PM@aOadbN6@qr@hoy3uQh6<O8\\\"\\\","));
$write("%s",("2):f(\\\"\\\"{ZpQx*opxz9Ps/3c:a4XYp=aUzTq;*e\\\"\\\",2):f(\\\"\\\"{u,M?ubFaF/gvdb|b8uJh>vgJKSm?6b7bM9Pa\\\"\\\",2):f(\\\"\\\"{vg(Dd#c/d4NuKL,@t/y,vE\\\"\\\",2):f(\\\"\\\"}Qa*bwbINZzxLUB3:tLbF1J+bV7-hTp1Y9v8\\\"\\\",2):f(\\\"\\\"{JnprZa=aIhBx.\\\"\\\",2):f(\\\"\\\"{X5/QPMWqz0;\\\"\\\",2):f(\\\"\\\"}Fqhb1bz0;\\\"\\\",2):f(\\\"\\\"}?NIZdtSaTF.dTa3y;<Bq.b3P3w?aY2cbG/Io49/byr.SWad0ebWa+eS\\\"\\\",2):f(\\\"\\\"{Ba9bP0TrjbdKpX+b9bt,6b>;Zw/bt,@QE\\\"\\\",2):f(\\\"\\\"}SaTFib.bpCgqSGSG.y6Web\\\"\\\",2):f(\\\"\\\"{6D9>Fa^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'aMNeX3s1\\\"\\\",2):f(\\\"\\\"{vft4MsUaUwC4Ga.SeXWxX7,Sf:~Xa*a,b?a:JSLtfbb3q;*Wau@bbA-:-\\\"\\\",2):f(\\\"\\\"{v\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"{LI7?ISa\\\"\\\",2):f(\\\"\\\"}~NftaXa0zXX|btvbb6b^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2):f(\\\"\\\"{#v3mja51(f\\\"\\\",2):f(\\\"\\\"{#,4353(za199(f\\\"\\\",2):f(\\\"\\\"{#(ntnirpn\\\"\\\",2):f(\\\"\\\"})215(f\\\"\\\",2):f(\\\"\\\"{#)|4[|4anb\\\"\\\",2):f(\\\"\\\"}s\\\"\\\",2):f(\\\"\\\"{yVRpRW*qNcEQxBa:.tv6wC4GaDQop<aD3bb:JabK:JQI|1j@uXuvvrB\\\"\\\",2):f(\\\"\\\"}wOhW-Ew45?9<abEC-mb?9<aFa8zvwHrV|h6vv>v>u7UaHazCoxTaTF/bKxdwW*ZQ\\\"\\\",2):f(\\\"\\\"}p,936N,JH>iQaBy*-iv,\\\"\\\",2):f(\\\"\\\"{7b5pyuBFwb<>urbv\\\"\\\",2):f(\\\"\\\"}r@W59i>59jg3b[aEG@f+0StS4-bf=jB@:5zWn>w<wrk\\\"\\\",2):f(\\\"\\\"{yzbXauupy?|6wfu186u1bi/Wa9bSaJd-KYzDo1jiRQlcb7Nh.*AAa2Ym:H8ezdZ001M4t<duwtgbu;1bEah,NJRaJd4JGaXRhqfb7qxjeLjy?o+5>;Z0Ps1GZ?Sr|T?ovpzzO0BVmzoRwby7VaV7q<ubD6n<:MvbfbrkK;H>RaVaOaM=mbe"));
$write("%s",("u:\\\"\\\",2):f(\\\"\\\"{SHxwt1fWa1F/Hp?\\\"\\\",2):f(\\\"\\\"}8;WaEaSyRa7b4-qs|TV\\\"\\\",2):f(\\\"\\\"{aOfbm?j<|btp42+F96fRtoGX8wu1hlp4bumbbY3.QawItp42WZEaRL1L1Xr/+F+b;rYakiy-TxpzEatbFaCYSpv55.w.QaBX5EFai>tW.G5>tKL21XDa*-NaJZfRL5lbn-&6eva.5Ba-bvAdbWiOGybmOgb@xXr^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'a@a4b8bc\\\"\\\",2):f(\\\"\\\"{>,A0Sab<ybRa7+Wa>a2;|-hb-so3a&aw5vs9+O08>,t>aq?cXT+4b\\\"\\\",2):f(\\\"\\\"{?<aB7W4fbOj6b9aB17Ah?L>jo@|6o-PUaWabr>a1tyWX|Fatc3b1v2;M|+6y?N1As6.C3c$bTa+GH>c9n5B1?a=aU|W|UaE2-s>atb*bFHxjEao?1;VaW>kiLV=?3bHZM|Wa9bW,hb-s:vs16JO0mb1<+F;v2-WaAaF|hboAI9rO8oAx+:EaTy=11VsJ+F66eqd8N@75/1X3VF7+bl"));
$write("%s",("wZ0OCtQ*b=Eq<ax|bG2kihOCYa8ub1Xgbo3F9\\\"\\\",2):f(\\\"\\\"{O1Cy-ubuAZ*yArg=qmuv3Dp<aOamu6AB*UnVx0bq<A*ZA|@2AM@3H<tg<L1\\\"\\\",2):f(\\\"\\\"{byX2..J*Le\\\"\\\",2):f(\\\"\\\"}Oto*wbhr42Eatb\\\"\\\",2):f(\\\"\\\"{6/+I2tbk3Eahx:fjY>xZ0Xa5G172Y*Smbg1mbxQ5.w.D45bkrtobbt/Pcdw*.LqbEQtNqLQOtdP0.3-oz3J\\\"\\\",2):f(\\\"\\\"{-R;RaAa1M6X/YK;Dvq?|-TaWa*3=a6Jv|Oa8o0B/@IoqC:6:\\\"\\\",2):f(\\\"\\\"{?ae\\\"\\\",2):f(\\\"\\\"{0x6d;aI72QU8VapokbBUpIXaSaR?vb8<Iqa.y,RTM*y-vXJxYg/T+dWaybAa|4c9c.EU=|5028o.bvqIQPtdwzPIoYa>ul;xSzb>\\\"\\\",2):f(\\\"\\\"{L|IK,b0bs<Zzpk/b/b6*DxYsbbn:@oVR@|mb5.\\\"\\\",2):f(\\\"\\\"}5VpPN3bX:,tI\\\"\\\",2):f(\\\"\\\"}j-<5lVlb9\\\"\\\",2):f(\\\"\\\"{TaAa3VcJ6bq<kihyj4K2swW2ERI\\\"\\\",2):f(\\\"\\\"}v50g1Tq7=s;s9s,\\\"\\\",2):f(\\\"\\\"{AsVPVa1YGrUa+dyFbb7bIq+bN|-b:Z>rjBcSG\\\"\\\",2):f(\\\"\\\"}X3.6m<B3i>3rPU*;|uJ8Za7bVnJZ3bs93bytvD4|P+ki/3A9eyaVa|bsqUDA-1\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"{|r*5.+Gv3bDyC3a7a9b2bBaPUDvfbdb>akbK3@QDkW6;vz9e\\\"\\\",2):f(\\\"\\\"{Yn+bAqv0oUD+Ea/S/3S3aSa<?e6-bOa1s1\\\"\\\",2):f(\\\"\\\"{Ec8\\\"\\\",2):f(\\\"\\\"{TXeV@azzL9cM5bBxY6m@|bHNbX<Oe+opOT*9@C5p.bRvw/vs+eF4F.;:JKCYdbnJaQaEpIA?+ZaZ?L<:Q:.-Z9v7L>GLII4SLdH-bub\\\"\\\",2):f(\\\"\\\"{E6/,b?+Bx95OaAroAjbeq/vLII4zvfbK2Cagbld5Ec\\\"\\\",2):f(\\\"\\\"{a?.tb,H>zo|:p6,OHlJGLTaPOPBsMc[a7PKLI\\\"\\\",2):f(\\\"\\\"}pCn5T\\\"\\\",2):f(\\\"\\\"{6u\\\"\\\",2):f(\\\"\\\"}+H9abby/va//-+yWvbb-bWa=\\\"\\\",2):f(\\\"\\\"{V\\\"\\\",2):f(\\\"\\\"{As6b70SaS\\\"\\\",2):f(\\\"\\\"{TFlbYHD3bbQa,4AaT+ibLZ5Z0|nx@UtNd4fDggcd?wBm@Aq=:iH,;GrNL+0TaOty?tsu,8oBtkrV2gF2Hy7Var<p<V\\\"\\\",2):f(\\\"\\\"{WnyblUVDbbmuvbF/>y*wAaAa7\\\"\\\",2):f(\\\"\\\"{-P\\\"\\\",2):f(\\\"\\\"{z+:mbyWq3FGqNEEI3kr*EFH96WZ3bn@gqYn+wxbYa8\\\"\\\",2):f(\\\"\\\"{tbG\\\"\\\",2):f(\\\"\\\"}cSD.h0tbYgMzBzyPSGZai9CEMqzr?|@aI|dHq*fGP"));
$write("%s",("aU8CEkbM18@99eRbCa<aXxdbxIbbf3-AufabIw,b@ozb*wcblbBODkwG<aEw4tE*mJwGF46-ID\\\"\\\",2):f(\\\"\\\"{LCaDvfbCafz8oT@.bN;.K*w?Ec\\\"\\\",2):f(\\\"\\\"{JdM.2uE*R>cb4berfbBafz=IYxSaT@/H3bR>cblbEwM2B1fbBaIKX1E*b3:sbb7b9\\\"\\\",2):f(\\\"\\\"}X1dZX1\\\"\\\",2):f(\\\"\\\"}scbSc84aIa8LuzQxUamIR>cb:6wGgJ\\\"\\\",2):f(\\\"\\\"{L0/,4|b.KSaGIab8oGIabki/3AaoGK|+2vbn-PaqNOa.F/Dc3s+awbrA2uki*Wh5wx3y||\\\"\\\",2):f(\\\"\\\"{b?Ik\\\"\\\",2):f(\\\"\\\"{Zav<EaSGZN/=:R26c0dd0im:*|s-FSymPub-=GvlbGibb\\\"\\\",2):f(\\\"\\\"}.ubcvVa@?ZqD9h*GvqzyT+elCvb\\\"\\\",2):f(\\\"\\\"{bZulb*;OTAqkiBl\\\"\\\",2):f(\\\"\\\"{bZpNazzG/Bxy9\\\"\\\",2):f(\\\"\\\"}odbOw@oWx,bXa/r1b=a4bkbubrAN|ub=w0Dr+hbcb3I3\\\"\\\",2):f(\\\"\\\"}0yw0KnStK|GvmbVwiICa?avbVPpS9N1bCaPQ.0GaDQj@I9mbpLjW>anCOA1GAIGvzbPa1jf<:iXQA8Zuv=Vwl>-EXatburAyM4Na@:tF1vG/Bxn\\\"\\\",2):f(\\\"\\\"{Nx-HvQt404QawIly5NebFaohVCBaU\\\"\\\",2):f(\\"));
$write("%s",("\"\\\"{jY>aVCb1F.8b7bcbbbAa<aMFX3Ua4</bl:eKaYazJ>p2bVa8ofb1LDSeq5/5:J8ybybmbHJFax>Pz9\\\"\\\",2):f(\\\"\\\"{P*BaPp?tDvIQUYcb<aiI\\\"\\\",2):f(\\\"\\\"{yZaXJ:;%3eKa3<+b2b\\\"\\\",2):f(\\\"\\\"}7K0Aaxbk5Njy-2b|TE0B|s2\\\"\\\",2):f(\\\"\\\"}udwPFpzjK5yNZ?rXaCsF0Va8oO4I>sqabLIRp>SjLaY2t<Va-xYl-x4b6-X;KEZzZ|1GPQyujb@C6F@,8TAr\\\"\\\",2):f(\\\"\\\"}IwbcWbbEa3bQ|.ykrpLHJc<24OadPrq0B@1<s:sOj<a|bm\\\"\\\",2):f(\\\"\\\"}LB7WTa3HvrNsI<bYRa/u5/-p5N6LloUJ=F52x\\\"\\\",2):f(\\\"\\\"{6@:VS5*X|bpVnN-ylV@Ukb*b0VpOzbFazCYzYaO/TqCIh*-.gWqifbgb@,kb71gf<.<OzuTrW*>we++bk:CK.1K,42wb=Rd|dzo;nC\\\"\\\",2):f(\\\"\\\"}sxb8bko>M\\\"\\\",2):f(\\\"\\\"{tttjbh2K|zbgbUaBaiON*YFG56gq/iO3<9-ixXXxbPqcqx+*bH=MmF+|lYXWXab+RubZafB8:I\\\"\\\",2):f(\\\"\\\"}4bZqhDfDzbPX,z5.cbxzXwmb-7+ThvF+CauT1;aye-*4EXH=Y33bFax+0yU*\\\"\\\",2):f(\\\"\\\"}b+b34H=RLVaxbTw3VTy615syb.bWaNqh*gb2.\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"}+.<P5?T.<=TmbMnk\\\"\\\",2):f(\\\"\\\"{irgDHx/pPaRT9y.yvbXQNa>7wb?oE*CwDvIrDvV=/b3PGa3CkbYx-bgbfWRW<WOW1q?*HsKxDxx+NVyrO=VD1|xA|9YnS3,\\\"\\\",2):f(\\\"\\\"{F/P9vss68bu4b3NaB*U*-9Wns6cbDvv0\\\"\\\",2):f(\\\"\\\"}B0BWaIri=\\\"\\\",2):f(\\\"\\\"{I5OfhAanxecmNUD1tcbtbhwMoBBez8ox+UwibINecqrzK?:\\\"\\\",2):f(\\\"\\\"}b6b9boRVwldUDF+UzpFyvC.mu8z6zLo2wev.x8zlt4zVwd5Jxhb8Tv4opGaL**JasPpxtOaLzBuubfviv5lU5BJ>TAL>B9PjcFaPafbeb+b7b6LX31sybVaw@5/PF7vVw\\\"\\\",2):f(\\\"\\\"{6k\\\"\\\",2):f(\\\"\\\"{fvt2?\\\"\\\",2):f(\\\"\\\"}HzebArdy04XKqqub9APadbJqt80b|b,bUq8871\\\"\\\",2):f(\\\"\\\"}zbEozt3q<N2p4dbhxpO+bs2PPQa*u\\\"\\\",2):f(\\\"\\\"}/PFXqy6lE6FGiFHDi>aGaoSJ8y7Zr:\\\"\\\",2):f(\\\"\\\"{649I/sFa>a4<sUi:,q5b-56b\\\"\\\",2):f(\\\"\\\"}ClQSTW7zPmH+xTB=\\\"\\\",2):f(\\\"\\\"{qN2ttq=?Y-i=bbX?F0jzib2b/rXSlb00;qOAXF*bDqmb1AdbrysJiRt4+9<>L7Jx96Ua@aC6y65b\\\"\\\",2):f(\\\"\\\"}"));
$write("%s",("pI:to0HfR@aHv409fxrab8@zqS.935@S.7Rt2eb=a-bXa1P-s+cqRt>|b8oZabbq*YtFjF2Ho3pjbW2<afbi|\\\"\\\",2):f(\\\"\\\"{bGxmbD@sszx-A+xZaL|,r-w.FLry?ldkAmShbjbtqzzZaBSkb@avsv<U6qNDr9b1b0-?f,8m<Yh8o|z?*nsQ@9b0bgvNa|b43Fy32Sa9bxrluw;2b8bYaIQ4bdb6bX>cqu1ki\\\"\\\",2):f(\\\"\\\"}RiSuwA5hbXaOwTaZs@IOa/kI8mGaiSvK2mbki6IiO\\\"\\\",2):f(\\\"\\\"{bSt8=PskiqG2|42tbb7yb9bRvbqi8w=\\\"\\\",2):f(\\\"\\\"{uBa\\\"\\\",2):f(\\\"\\\"{b**Zq8bC:tBybZzFHPaOa5bY?Rn5b7pb7IQCx1<lb0vmbe\\\"\\\",2):f(\\\"\\\"}vbFjgF.<;DBL8POao-e-P6-7NCV4k4E761F2F+iO2bFri9ZneJXiWa?a3b3,+c0bAa*b3bHMc\\\"\\\",2):f(\\\"\\\"{1bvr.bzblI3bjbb*dkPalQ-2wb\\\"\\\",2):f(\\\"\\\"{uQa>v5E*bbuLQV4Nafb01EPu44b-jNaPaYh|pimkil*?v95ViZa2Q<a*EC-,h*bpOwbz@0N2b5\\\"\\\",2):f(\\\"\\\"}YIBaT2ZaSa0NNw5EFF*b\\\"\\\",2):f(\\\"\\\"{6or7\\\"\\\",2):f(\\\"\\\"}9y9bdb|s6bNa0bS=VnIuQPxjTa?\\\"\\\",2):f(\\\"\\\"}+bZN1jIpS0v<7\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{d9bAqGaGO\\\"\\\",2):f(\\\"\\\"{u;qG.;tvb|sN6h2L9v<Sa\\\"\\\",2):f(\\\"\\\"}bUa\\\"\\\",2):f(\\\"\\\"}G\\\"\\\",2):f(\\\"\\\"{JNabb>r,bkb</s2Aas7ib</kb+4ItCpcbOu=3?L;NNaI4Xv5nfb6zxbdPbov|mb?awzK431Z,c2TaFa8Nu4C0DoL\\\"\\\",2):f(\\\"\\\"{/1fhtb7b\\\"\\\",2):f(\\\"\\\"}L::m?41=aXxQxybgbAyTxfb0b-KK@2bNx8@+bRB5,f<\\\"\\\",2):f(\\\"\\\"}oVmWqYa|5+6ab+b8bS0sqkiJu8O6b|b0yyF31XxJnkb5,mb@o1GVC\\\"\\\",2):f(\\\"\\\"{Ohtk51x9bN|Zwi|B\\\"\\\",2):f(\\\"\\\"{*byb:-x+/bp|hbWwXaHI1bA0Panr96N1TaV+irQaZa+9gbdgT>Lq8oUaOANnc;G\\\"\\\",2):f(\\\"\\\"{wbOavbQaTaOl|bzdW2d/ZaPaPzk5wbnKjb*;PaA<a>Tp,bgmuqW2HtXaMhV:PakGub=H?J8oVa0b/b,rhb7bjb5/4z-bAK1q/q1b17hqYt<kx3ybe41;tb0yr*Ir4b9o/GEpY6u1+6Cx/rDaX4P8jbR8P8wz4pV;0pTp@,>,bbPa5.-bTaCxB*\\\"\\\",2):f(\\\"\\\"{bXa-\\\"\\\",2):f(\\\"\\\"}4e.xM4o+jbA<D8Xyf\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{5-rosjI*23o8b./>a<aV|gb1oS"));
$write("%s",("wF4=\\\"\\\",2):f(\\\"\\\"{|oTaeM@a<>uo-bNsAvDCn-4bYiJkKtCaQoxhy+eb<al0=ay2VI/I9bAa<>yJ7uzv|r@@V0+bUimbfGgqoudbio+\\\"\\\",2):f(\\\"\\\"}-=/5-5-pwb?3Pzq?yb=|8vDazbDy*tjJ6s.<CJ=B,<\\\"\\\",2):f(\\\"\\\"{:V\\\"\\\",2):f(\\\"\\\"}/>v15zXqOrMqcbUr\\\"\\\",2):f(\\\"\\\"{bjbI\\\"\\\",2):f(\\\"\\\"{Ta-b7bmbXawwpxY0\\\"\\\",2):f(\\\"\\\"}bxb=a1brsQabbqIvbzCF9f0Ms3hlbI/Xap+*>@?u49gWrk\\\"\\\",2):f(\\\"\\\"{8CQaEEZa:6VCJz3oEyuq+bkoltai-b@+ax-iJ8i1yFK|6b::mbYa9bHgc+l:\\\"\\\",2):f(\\\"\\\"}=XxXr8o*t96S</p>,:suyJdu;3IdbQ/jl|bSyd,Q6D3ubab-bwu@Iu:t*7b0bhof9D3SG?ayb?axt;pxwF\\\"\\\",2):f(\\\"\\\"{8oh9<a*wT*M0cbR@kbPJ?aGasxeq\\\"\\\",2):f(\\\"\\\"{y*zC9OaabMq<a@akiD/+b,|8bz0AoWpOjebtbom4b30S.|1-</l9D=H7bmoBD1\\\"\\\",2):f(\\\"\\\"{2bo\\\"\\\",2):f(\\\"\\\"}/bt<@aq/mb.b5;/b\\\"\\\",2):f(\\\"\\\"{or2/bEafz4.|b.uF/,\\\"\\\",2):f(\\\"\\\"{;qAa-bZ|yFub+bOaq.Y8tAfbyw\\\"\\\",2):f(\\\"\\\"}|mr\\\"\\\",2):f("));
$write("%s",("\\\"\\\"}tKHMq2p.b=qNacH8o\\\"\\\",2):f(\\\"\\\"{E7B\\\"\\\",2):f(\\\"\\\"{bNa/*zbEaPaVa-z5>CyiFYaBo|B0bD5Ua|*fb?awbm\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{sVa?\\\"\\\",2):f(\\\"\\\"}Cx0bFa=1CalbYEA0Na;sHo8beBb:*b1pCnlC|bZ4X4M64bQxjbKtjbXs.p>a1bf5qibb+bwbQaFaADQa3bs>OCabRaM1Pz?Dtbqz*>Ktezx+Urm@ou>qCxaGgb2bvboxb3/p*t>w?aA17HQxTaRawx\\\"\\\",2):f(\\\"\\\"{bOargIoI7u/4a;Hgn;FDtcbDGRaBfEFJ=ybd4cb.bSaqCDa\\\"\\\",2):f(\\\"\\\"}b*.Paf83p:,pzaBc.43KF8vHgx6095bybdb2q9b<aUaODDaVaU9u4|@hbA<RxX\\\"\\\",2):f(\\\"\\\"{XB5tE.8GC:kb|@*bnqu-<q>aZ>/sgbUrwx>9ybar\\\"\\\",2):f(\\\"\\\"}b.b,1H>?0Wacbs1U9dAa/\\\"\\\",2):f(\\\"\\\"}-E:f:VaZa|bvbAaXaIDFakib46FTa?+RaB|\\\"\\\",2):f(\\\"\\\"{b*+Wv-b0ba0Qa@a1;K|S@pC>a.bjb8oubyFloCrn3qi|5zb+0Pt82*93b\\\"\\\",2):f(\\\"\\\"}bgb|b2\\\"\\\",2):f(\\\"\\\"{uxNhPaw/Fa7>8oRa.FFa8v4<?h=aDqz/Ta=EAy17VaHwr,f8K\\\"\\\",2):f(\\\"\\\"}Va-l9Fdp7Dv0A<YaG"));
$write("%s",("ajAm2\\\"\\\",2):f(\\\"\\\"}tX\\\"\\\",2):f(\\\"\\\"{uzvFlb4bv0jbw5Y,Y?i9Bacbq-Bav2CpRa\\\"\\\",2):f(\\\"\\\"{6kr<a/b5uxtFac.8b=A<aO|-bUahvK.gtBaTBjbI7-AC.gbv0*\\\"\\\",2):f(\\\"\\\"{Cw0bg1SaPt*zj0Ba8=9bh0i=g,h*xbe6>ag,5gxt1b5uybzbg1j38@,o-dAvybw/z6OaVivpa.-bFaEpq*|bWvL,@a0bfb2gI|GrXawbQz0bOtkre+IgYu\\\"\\\",2):f(\\\"\\\"{be<stA*0zdbGrCr3\\\"\\\",2):f(\\\"\\\"}@|7b3hy+F4b2+bTafbWnFz,2k\\\"\\\",2):f(\\\"\\\"}y36b/+ogFyIoNC/b/zI5*3dbY?dyOaAaOz@a6g*2S.\\\"\\\",2):f(\\\"\\\"}:v\\\"\\\",2):f(\\\"\\\"{;B5l9Byw0bm?n9Ff|3PaCaO2bBe9suUr4,;vO17A;7BBq9+Bm:zvH=qvibEa8v<\\\"\\\",2):f(\\\"\\\"}4,Xal\\\"\\\",2):f(\\\"\\\"{WxibbubbC+w+?,kb1b/*\\\"\\\",2):f(\\\"\\\"}|X*ebvqgbP;,b71Wy8;m3ab|bFBkiOo/COaQyK3.b4p@aXsgf186bBfY:pCJz-rf:hh.bR;Wz=aI8BrwxkikBiBouWaL|V0Ea?\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"abyfr,b\\\"\\\",2):f(\\\"\\\"{9Twzuqu*bcvZ9Qatb8o-\\\"\\\",2):f(\\\"\\\"}5bav=atoNvebbb3s<8x5v5kbAtZui;"));
$write("%s",("/sDa/*7A9pybWatbjuybxbm\\\"\\\",2):f(\\\"\\\"}Qaj00y18/8-8+86bvpY8\\\"\\\",2):f(\\\"\\\"}b7b?qc+in.<<3T\\\"\\\",2):f(\\\"\\\"}3@2l1@V;9bFah6.b@pP9Ta0bQ6I4ytwtutstytQ/Y3qslqQa=a2-ib=a5bSa3\\\"\\\",2):f(\\\"\\\"}=wzdLpb.Euj6Yahzrkgq3bXay+\\\"\\\",2):f(\\\"\\\"{bogXaUaubA<=a6\\\"\\\",2):f(\\\"\\\"}*b>a6\\\"\\\",2):f(\\\"\\\"},xTaz,Da.+9b@thtz@i9p+A*ZargwrJxd5-9r+Zp|*-by+Z*z,hbmu3b@ak\\\"\\\",2):f(\\\"\\\"{+b6bTpxb*Y29-.u0Nad5h2\\\"\\\",2):f(\\\"\\\"}bvbG3om-9r,muimu1-b8bgbbbOa1bXa\\\"\\\",2):f(\\\"\\\"{bZxV7kiY7Io-bdbmuZwWa=*;<Z0D*l+*bfbP6*4abNa@iPaDk6,Pajt?oWyCwA8Yagq:-bv1b1qnswy2btrD3a\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{bb\\\"\\\",2):f(\\\"\\\"{.8z@fbOux1T55lR5.<->/sUa+\\\"\\\",2):f(\\\"\\\"{Q*fh1bj>D1-bDa-bAfBazbjv3b>aI7abG5xzj0mbTaax@?Dapz>aYaF96*DaW3p->pbbYa<a1btbg=krbbWa03@,Syfg<aO\\\"\\\",2):f(\\\"\\\"{F4B95b1qI/Q39<,vDa\\\"\\\",2):f(\\\"\\\"{b-dwb-dW9>a2b.1+y:f.t3|D"));
$write("%s",("5G6Wa.bS0Asc,1\\\"\\\",2):f(\\\"\\\"{-r@<Dwb+hb4ba.+6hbEaf7n|tzxbm/,tgkAay7Ua3bCaN;yu>,VmX;K2V4N<Vab<8oWa8bN-?a1;mb@h|xK|@avb8otb59zbvb>aupSaWaD7|rvbSqez>a6>hw?aZr@7Faub24>a=a3bWo8bYqd5K2Ou5x|:n8*<5bW4A89\\\"\\\",2):f(\\\"\\\"{2*BaL9v>lbPa@hJ/Aa=ss6x:Zx\\\"\\\",2):f(\\\"\\\"}bm\\\"\\\",2):f(\\\"\\\"}?a1bKpxbvb\\\"\\\",2):f(\\\"\\\"}b5/*bFaky?h|babtbk=PzNnjblbsq6b/*q7drU,CnFau\\\"\\\",2):f(\\\"\\\"}m6-iBwOaduaqh=*\\\"\\\",2):f(\\\"\\\"{holv4|Xqgv;rHomrqqZaOaRa3powz,5bxwVaf+iwDao\\\"\\\",2):f(\\\"\\\"}hbD41*/*-*|x-*Y+v=+plbEa?,?02|\\\"\\\",2):f(\\\"\\\"{bF8A<>7\\\"\\\",2):f(\\\"\\\"{y*bXa8o88,bJ\\\"\\\",2):f(\\\"\\\"{|bmbJn04Dp<:FxJdxr8b=pOa@pJv\\\"\\\",2):f(\\\"\\\"{bV0u\\\"\\\",2):f(\\\"\\\"}uzVa@aibcb1tCx,b2\\\"\\\",2):f(\\\"\\\"{:vAqIrk|J\\\"\\\",2):f(\\\"\\\"{TpTa\\\"\\\",2):f(\\\"\\\"}5Z|Wa-9Gs-bG2+dDa8bo;t.2bEaCwTa.<m8X.R.z1:3z:\\\"\\\",2):f(\\\"\\\"{b+5u,/b@,XyomkbUtWa0bJ,?a9sRpTpVa"));
$write("%s",("*+*bhbt1l\\\"\\\",2):f(\\\"\\\"{2bCa7|>t-t<ai/,ha.EaI-,birB1MmWa0*mbW,8bl.VaWaSa\\\"\\\",2):f(\\\"\\\"{.O\\\"\\\",2):f(\\\"\\\"{S-o\\\"\\\",2):f(\\\"\\\"}Sp2+V\\\"\\\",2):f(\\\"\\\"{E7\\\"\\\",2):f(\\\"\\\"{b*3K-ebB1Ta=\\\"\\\",2):f(\\\"\\\"}59rqUa?q*3*;Wa=t3bubHtbr|;Aa.bQ+abE7VaF7I-F|t1@aV7\\\"\\\",2):f(\\\"\\\"{blbIs<tkvaz1b>a\\\"\\\",2):f(\\\"\\\"}bSaPz-\\\"\\\",2):f(\\\"\\\"}ybhwT\\\"\\\",2):f(\\\"\\\"{,d\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}y\\\"\\\",2):f(\\\"\\\"}tb7:l6B3.0.bxbZh18FxV38\\\"\\\",2):f(\\\"\\\"{XxHpyx,bCae9ub62wb.rqrQaVaPxzbB*w,Ua.b8\\\"\\\",2):f(\\\"\\\"{;*7bPy*bE6eb7b+8OtwbSahhu6,4H\\\"\\\",2):f(\\\"\\\"{Wwwt;5?ax\\\"\\\",2):f(\\\"\\\"{Su;3-,o8,tfb@aYatbFya0Xya58//w7bOaD|.*p-G-/w6zAaCtG\\\"\\\",2):f(\\\"\\\"}jv\\\"\\\",2):f(\\\"\\\"{bpx@a0\\\"\\\",2):f(\\\"\\\"{Af,bNnebktX5h0,5fb\\\"\\\",2):f(\\\"\\\"}b<83*lbBqY5fbFaGgwb=vablbWaCaP6Aa,b\\\"\\\",2):f(\\\"\\\"}p>ahw3+tb+bmbkrFa/bo/Sv\\\"\\\",2):f(\\\"\\\"}bjbQso/Oay"));
$write("%s",("bZakb@,lb?aPa-b9z023|Mo/pt8/pxtvttt+b2z|b+\\\"\\\",2):f(\\\"\\\"}Ga@23\\\"\\\",2):f(\\\"\\\"}-\\\"\\\",2):f(\\\"\\\"}H\\\"\\\",2):f(\\\"\\\"{5b3bE7.3E-omxbHuDvFavbW|UoXvlbDaBaTahzPt8\\\"\\\",2):f(\\\"\\\"{/bkim0?+tb5|+3DaXq\\\"\\\",2):f(\\\"\\\"{bvsE6ibmbxbZ\\\"\\\",2):f(\\\"\\\"{eqDaibwbFa?oG\\\"\\\",2):f(\\\"\\\"}k*o5zb5bOa*b|b-bSaK,cb@*q*\\\"\\\",2):f(\\\"\\\"}.8o/bT*T7ub\\\"\\\",2):f(\\\"\\\"}bVihbZainl8Q5T.O51\\\"\\\",2):f(\\\"\\\"{BakiB5P\\\"\\\",2):f(\\\"\\\"{Fazdyblu8zZaHoBaGaH*Zat|A-Kfib+bYna.7b\\\"\\\",2):f(\\\"\\\"}*DaZpfu\\\"\\\",2):f(\\\"\\\"{bfb*4VaTaTamyPygqkbyteb,bzoubRa1o/b|b?um6k6FaNa,bVm>u.61b8bt*l7KvL|*6Gag7D-O4J|e-Nakbl74bn|1bDao+Ua9fL|Syki|6Ra@aLnZ4abl6a\\\"\\\",2):f(\\\"\\\"{|bebY+5bWyOt3,3zcbkb:.hb,bcyFnh5z+QaYax|ub|bib=-Hd<5Uajtk*evlbwbRaB*6b8bf+@hPzw6Vw-wmuwb*yh5mb9b8ovbzb>aFaQaOaY\\\"\\\",2):f(\\\"\\\"}3bjumbix3bdb?u9blb7bibab8b2bkyWxhbqr3u2qlbozZa4bH.2l"));
$write("%s",("W.\\\"\\\",2):f(\\\"\\\"{12lR\\\"\\\",2):f(\\\"\\\"}S.P\\\"\\\",2):f(\\\"\\\"}83lbdb4bPz:uyb0b7bQaVwEa8ogbeb>apo3wqz9bcbF\\\"\\\",2):f(\\\"\\\"{-bn2Vazqq5Yao5/pl5fzqodb9-jb\\\"\\\",2):f(\\\"\\\"{bcb\\\"\\\",2):f(\\\"\\\"{b,bAaXxfb>aRaabxu@t5bg+x-|uVa3bXslbAaezT/8bE\\\"\\\",2):f(\\\"\\\"}Ba|f@ad4nh/b>a5b>avbDa=abvCaF3Sa>u7bpkfb@pu4Bo4bQc7b2bF/7b\\\"\\\",2):f(\\\"\\\"}btbF+.bh*Zxa0gb\\\"\\\",2):f(\\\"\\\"{4=|cxub+w+bvkJzabOaH\\\"\\\",2):f(\\\"\\\"{8bv.5bXaTaCa3b/b8gPaTa,bDaMombjbcb*/Ep:rubbchj*\\\"\\\",2):f(\\\"\\\"}4-@..bq.YrQa8bzb2b8o|bubEaebibi|gb?\\\"\\\",2):f(\\\"\\\"}1q*b-dybS2=pN*bbJn,bN2\\\"\\\",2):f(\\\"\\\"}bK2eb2b:2lbG\\\"\\\",2):f(\\\"\\\"}>aYtgfk*inS.w\\\"\\\",2):f(\\\"\\\"{Q.U.,,w1a\\\"\\\",2):f(\\\"\\\"{e3x2jbYq3bq+8oCaWa\\\"\\\",2):f(\\\"\\\"}b*b.bVaE05b8o3bNadbhtdb9y|bKxW\\\"\\\",2):f(\\\"\\\"{db1bebiu,bGaD\\\"\\\",2):f(\\\"\\\"{<a\\\"\\\",2):f(\\\"\\\"}+c\\\"\\\",2):f(\\\"\\\"}IdzbH23+T\\\"\\\",2):f(\\\"\\\"{zb/"));
$write("%s",("bf2L\\\"\\\",2):f(\\\"\\\"{1vyblboq4b*b0b>2+bkbQa9bzbDat*Oa50|bNahb5bpjvtkiDu=p2b7b3r/k;imb;r3eroFaTaWpfq=p7bhhvbkbtblbmb0\\\"\\\",2):f(\\\"\\\"{Lps.1bL,bc<|wbu1*b2bTaNa:|LhEacbCavbDnoqzb-0fb9b0rvb-bGrl\\\"\\\",2):f(\\\"\\\"{:1zbA|\\\"\\\",2):f(\\\"\\\"}bB/ezNvryioWazb4b@at|\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"{-Naevfb8ywbB*acUa5btbF|ZzNaPzB*4wYra\\\"\\\",2):f(\\\"\\\"{Fajb2|\\\"\\\",2):f(\\\"\\\"}bEag|\\\"\\\",2):f(\\\"\\\"}.kb;y+bSv*bVmT/x\\\"\\\",2):f(\\\"\\\"{/,8xx\\\"\\\",2):f(\\\"\\\"{6x\\\"\\\",2):f(\\\"\\\"{iV.2bjb=aWa8oM.j1<aNa7+M.|bZaRa/bjb0bhb8o9btbXaFagblbA-gbK/KnNaFaEv=aFahz?a;t5b,j6z\\\"\\\",2):f(\\\"\\\"}bYa2b<akbYa@hYaeoAa@o1tf\\\"\\\",2):f(\\\"\\\"{?pjw.0NxSa,nfbXaXaPz?pabxt/bBav0hbwb=a.bTreb-b3uFawbZahb=aBaZaq.ibm*dbvbluCa3p?ax-tbsqvbmu-uXaSt3b2|Hn1bBvOa=\\\"\\\",2):f(\\\"\\\"{ib3b=pgbgwZaiuc\\\"\\\",2):f(\\\"\\\"{*b/b/*vb.b8o<a\\\"\\\",2):f(\\\"\\\"}b/bPzir5y|b"));
$write("%s",("U\\\"\\\",2):f(\\\"\\\"{Yairtc1|?aCa9b*bSaTxo/+e+b=aNajv2kzb*b+b,s.bub8q6q.bK,ab-wabUa>aL-?asoUaOavja/RaG.E.@.>.lb<.Sacb8oyi+,:x.,Q\\\"\\\",2):f(\\\"\\\"}y\\\"\\\",2):f(\\\"\\\"{O\\\"\\\",2):f(\\\"\\\"}U\\\"\\\",2):f(\\\"\\\"}7xucwb@u?aL-EyV\\\"\\\",2):f(\\\"\\\"{p..bBa@a\\\"\\\",2):f(\\\"\\\"{b+bRa/s=aSa=a/bE-Qa..xbCa4.=aab1bRa4bzb0bRaszez.b0bjb:v=aVau-Kteo<a3bBa>a\\\"\\\",2):f(\\\"\\\"{bibRacbDaS-<aWalbu|N\\\"\\\",2):f(\\\"\\\"{cbVaVaO,Ra.-wb/bVaPa>aEaAaOa=a1hRaxh:\\\"\\\",2):f(\\\"\\\"}=aEaezQlE-TaSa@agbNac\\\"\\\",2):f(\\\"\\\"{Ra.bmbybvbuy6->aSa0h\\\"\\\",2):f(\\\"\\\"{zXaabhjOalb@aWaWaTa<aEa.bRa/v@au-SaVaSaAaV,TaHnkw\\\"\\\",2):f(\\\"\\\"{|?aUrCo?oabubLn7bAaayib0bg\\\"\\\",2):f(\\\"\\\"}tpFgto0bibebCa-xPa.bSqSa8owb>a+bot\\\"\\\",2):f(\\\"\\\"{oot6b*bNn6bZa@awbBn/b,s6tFgtpRaFaxbgb5babd|ZaAa,t8yDygb0blbUa+vxhOu3l*,s\\\"\\\",2):f(\\\"\\\"{enS\\\"\\\",2):f(\\\"\\\"}N\\\"\\\",2):f(\\\"\\\"}z,lbs"));
$write("%s",("z+bWzA*,bTaOa2bUrNaU*Zp5bbkpzjbLy>xVaFa8ok\\\"\\\",2):f(\\\"\\\"{-i1berlbm*abbbUa1bVaub>a1vV\\\"\\\",2):f(\\\"\\\"{EaNa.+oqwr\\\"\\\",2):f(\\\"\\\"}w\\\"\\\",2):f(\\\"\\\"{w0z>x.bylhbbuBpUpldg*\\\"\\\",2):f(\\\"\\\"{bmbBaSa4bhbWaUa8bEa8bVa4bNaFtNr*bcbOahj\\\"\\\",2):f(\\\"\\\"{bSvCaebnwbuQa4bYaDaubWaxj0ydbbbkbCa,bPa?a2b+t<a6bXacbcb,b7bkbGsUacqlbkb+vZaUaB\\\"\\\",2):f(\\\"\\\"{lbmuRa2bOakiRw<a=akisr<aSaBa,b/|Oa,b*bjbOa3bSxPafhCa?|\\\"\\\",2):f(\\\"\\\"{bUazuBa6bnwTaXabb\\\"\\\",2):f(\\\"\\\"}babroRvVw0b6bZv0b+bjbUxLsebzbe\\\"\\\",2):f(\\\"\\\"{kbkbgcUoZt8oeb8b@ozpTa5bGgXx=a>tefybEaubItinx\\\"\\\",2):f(\\\"\\\"{jsbn9xt\\\"\\\",2):f(\\\"\\\"{x\\\"\\\",2):f(\\\"\\\"{r\\\"\\\",2):f(\\\"\\\"{u\\\"\\\",2):f(\\\"\\\"{p\\\"\\\",2):f(\\\"\\\"{bbim<acxwb7btbebcbvw1b+w+tFa4b,hmbeb?albYaybUaZa8ook<axwHxZsyb9pfb3bkbazok1t3b6bbb|b-rib6b\\\"\\\",2):f(\\\"\\\"}bSpex2pwbvbwb\\\"\\\",2):f(\\\"\\\"}bCa0bruBadb*bfzjb"));
$write("%s",(".bibHujb7bLv<a?aNa*b1bjb3bZamb4bCaNa8bAaUa8oFaZtlb>vcb1uNa?aFa*bpoQa7b3gcbJ\\\"\\\",2):f(\\\"\\\"{*o9bbtZ\\\"\\\",2):f(\\\"\\\"{EaEadbzbdbkbluIkIrTazb3bibSaCrzpBaUaRagy/b*bo|m|=a\\\"\\\",2):f(\\\"\\\"{bgb*bib@qzubbCaab?abbab*btbYsUawveb|bRaubcbEapoXa7blbQaCqz2/bJdib6fXadw.\\\"\\\",2):f(\\\"\\\"{kiGoWo1bwvbb0zCadb/usu-bwb\\\"\\\",2):f(\\\"\\\"{bdbVa=r*bEaYaQa0bXzkbUabb4b5bEv0q5bOuPuq\\\"\\\",2):f(\\\"\\\"{Nuis;xgsOulshs4xDp8ovpkbPauff\\\"\\\",2):f(\\\"\\\"{NajbPatbSalbtbPawbWa*b,bGzFazrLzWrBaFaibDatbNazr0b,b3b,nybrgkq,bvbbuGuwzFaoxwbPxZp4bRafb\\\"\\\",2):f(\\\"\\\"{bbbFa3bCo0bUaxbtb8b8bZaXa0bSa0bkbxlPa2btpbb=aOaXiebSaXa8y+bybjxibCxxbAalbgb,bydcbAa\\\"\\\",2):f(\\\"\\\"{bly/bub@wwtmbgb4bVacbabWo0bVa\\\"\\\",2):f(\\\"\\\"}ygb\\\"\\\",2):f(\\\"\\\"{yyyVa8bwbUa\\\"\\\",2):f(\\\"\\\"{b.bOa+y\\\"\\\",2):f(\\\"\\\"}y\\\"\\\",2):f(\\\"\\\"}bKh=xzbIwlbBaOaTa7bbbybbbgu+b>afbi"));
$write("%s",("bEwRakbVaWwibVaYa0h6b1x3bSatqTa3bWpvbSa/bDaybfbnxQaUaduxbFaYaeb\\\"\\\",2):f(\\\"\\\"}bmbubgbybOaQadbUa7bzbwb0bCa1xEx-b8o/r-bab\\\"\\\",2):f(\\\"\\\"}bNaYaZa6bBaxj5bBa1x\\\"\\\",2):f(\\\"\\\"{iipjpyihpOuQuOuRufbexgb/bAtPa*b8bjbht0oPaBtTaabIt0bebhc/omx6bPwdb0b8o*bvr0b8babxb7bAotbCa\\\"\\\",2):f(\\\"\\\"}b,tcb/babgbabFa2b1b8o+bNwSv6b,b8ozqkv;vXaNawwwbXaxw\\\"\\\",2):f(\\\"\\\"{b,jQr+bloYabblbibffYa8bhr*b;rRa5bfbPa|r5b1b<a8bSaCa8bxbEa0bcbFafb8oyb7b\\\"\\\",2):f(\\\"\\\"{bilUq/b7bxb4btbabcb8b\\\"\\\",2):f(\\\"\\\"{bebhlNq,bwt>pKrkbxbib>a8oxp?r5bZa1bIrzveb0btbjbab7bWqPakb/bUacbvbZa-pkb+bUactRa8bFaebab0bZsavZaivUaAaeb/bmbNazblb0b@t/bkbabfvBagb1j1bltFj5b|bVaetct,bdbRa1bkbcb7b.bur5b/b-bcb6bwb<r6b0qOuesMufs4aks1lcsdb8okb\\\"\\\",2):f(\\\"\\\"}bbbibzu8o,b\\\"\\\",2):f(\\\"\\\"{bWayubb1bfb,bHqQa\\\"\\\",2):f(\\\"\\\"{b*rdb,bWaxbdkEalbybwbEa1bWa"));
$write("%s",("|b0ovbYa+bZawbkb7bfbZajbecZa1jsploFaUaNaXago1b7bxj8bebXaDa2bmb6gmbwbLtZa<t8bbb0bctTa1bwb-j<aZrdb<tmbPahbgb\\\"\\\",2):f(\\\"\\\"{btplq7bXa-bkbTa@akb5brpQaxbNaVaQa?a+bvblb:ftbCo3bYa\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"}bOaOj?a/pcbmbEabbfbUaibJoPaEjRa3s0g8b0bubNa\\\"\\\",2):f(\\\"\\\"}bVatbfbcb5bjb0s\\\"\\\",2):f(\\\"\\\"}bTaZaCq,bFaogCaOaxbDaoqvb6bjb0r.rfbzb@a<rBq@qXaWaFa.b8b>idb/bSaubub5bNaxbVa5bhbxb@aXa|bjbRadb1r/rCakb9b*r|rzrxr@a/bPaubUawb@adb-binyifpdsgpkpepininMiYoZavb7bNaAakblb+bXa?ombCawq7b>a.d6bhbFa|b7bDa8ofhub8o\\\"\\\",2):f(\\\"\\\"}bDa6bdbwb5p=aYa4bSaabZqbdfg>aebnrLn-b\\\"\\\",2):f(\\\"\\\"{bubjb9b.b?aebAa2bUaGacrRatb\\\"\\\",2):f(\\\"\\\"{b8o0brqyb-jdbTa\\\"\\\",2):f(\\\"\\\"}b,bjb+c2bfb-b3bUaki-oValb\\\"\\\",2):f(\\\"\\\"{bwb2b0bQaybDa@a8oPaEaCoFa8b?a0b>aWahbZh\\\"\\\",2):f(\\\"\\\"}b1bdb8b.bTaQamb=aebQa|b\\\"\\\",2):f(\\\"\\\"{"));
$write("%s",("buqsq>aNalb5b@aFa+b3bDaFaYpWp1oYi5bEoyp6bcbMn\\\"\\\",2):f(\\\"\\\"{bkbdbab4bjbNaNhkbRaioubkbmozbebmbibTaDp,bOakbNacbYaabEajbjb|bhb*bBaDabbtccbPa,dmbAabb2bdbPabbDaDa3bAa0bdbAa>a,bcb>alb2bXavbvb5bcbOhTajbEaxb8oDakb=ajbtb|bEaZaFaAatb2b,bibOaXaib8o\\\"\\\",2):f(\\\"\\\"{iapbp-lZo-lcphn\\\"\\\",2):f(\\\"\\\"{ilnmn\\\"\\\",2):f(\\\"\\\"{ikninubPajbYavffbkbyb8oib+dbbbb,bebYa8o4bDaYadbYaXaBaabwb*bCaDaSnjbGa.o4oDahb+ogbvbNa1bkiqb7b<a>adb<alb,bYauovotoro7b/bYagbibjbDavb*bOaEavbdbFacbZa.b-beblbzb,bNa7bvbCaEahb<aCabb*b8hQaub*bWaQagbSa,bEa7b6bAaEaMl6nxn3nsn0nTmvm0n;aznwm?aumznAm?l*n-bMl8mCa>lQmwbic8a9m@lmmtnEaXlBmom>l|mjmhmin5l5lcn4afn9ayidn-lan0l\\\"\\\",2):f(\\\"\\\"{i4l/b\\\"\\\",2):f(\\\"\\\"{f-a;hub@hBm=a\\\"\\\",2):f(\\\"\\\"}mJm=l9aEaOaBm@m1m2i:a-bBmnh-a2m,mCaXlbm\\\"\\\",2):f(\\\"\\\"{m@a<a-b|e5m+mPllmamRlPlNlsm*m:aCa|exm"));
$write("%s",(">aAammWlRl9a;lSlAa;kIl|ekmxlMlZlBa-aOlHlFl*bvbtb/b-a+bIdAlTlBlKl@aIlMlSe|eGlLl?aAa>l\\\"\\\",2):f(\\\"\\\"{b<lClAlFa?l=l;lHa9l9a|e:lxb8a+e-a1beg8aXful8arb|eidxi2l2l.l3aLiyi,l-fzinlOhFf6b-a+czbxbubHaqb6aqbEiFiDi5aqb@g-a,bAfzb.bKfnbxb\\\"\\\",2):f(\\\"\\\"}ikiZgXg\\\"\\\",2):f(\\\"\\\"{gag\\\"\\\",2):f(\\\"\\\"}h7i@kvh>ktcBa3a;dLfbkAk4kWjBa?a3aPhIgDiwbJa8iDhZj*hXjDa?a>aKi6e;hrbckakik5jCaKi2b3bGiUfyj8f2iDj?a4jKa\\\"\\\",2):f(\\\"\\\"{b;a3gwbccIa3b1b-j,b|b0avh7hvhQiOiMi@aKiyb3bTj?a9j5i5h6jBaLiMf1i\\\"\\\",2):f(\\\"\\\"{g\\\"\\\",2):f(\\\"\\\"{gsbubwbki-aDjBj:a;b?j1b0b-b3aAa3a7b-aki.a:b:b,b7hWhPimiNi@a3a;hwb+b-aPcuj/b8b1bPcxb;aUf-b:fZapg|b.b5b-amj>i3bWfvb|bIgGipgfg3bgf;a<b:b3b-a8bIg,bxb2b2btb;a7h*h6iPa4i3a>a3a5anb-aEi/b3b4b.bHa8byb2b2gtbWfxb5b+bYg7h5hliYhWh;d+cKfHa-i-iFaGaji|fld4a.gwi/auh4a-afgdgMaFa=aWh-bYhDhChGa+"));
$write("%s",("bJdRh9a/b5a|fCc8g-bPaBaobDhHfMa9aMaIa5axb3b.b4b0bxbzb-btbeg7hkg5hGaMbHg2bzb;azbLfccJa7b?a?auh*hCdYaOaVafbVaibNa=avhvh?a;aSgVaNaUa.guhkgvbpbEa*c7b=aAaCaCa>anbJdubSczbPfIcQgyfwfuf2bsfNd3bHa?e-a-fZf:aIa+c9f:avbldub4bcb-b3ggc0gHaebdbJaGagfef8a1bxbwbtbxbUaac|b3bdgfb/akgzgtbxcRf?a1akg-a6a5bhg>azd:a,cNahgwb.b;b>aagob,c:a-a.b\\\"\\\",2):f(\\\"\\\"{bvbxb5a1aob,fCe2b-a:b1dtbHa6a/c2b/a,fPcFf/b:b6aKa6e1b4eIa8btb1b1bNaGatb5a+ctb,b-a\\\"\\\",2):f(\\\"\\\"{fyb3dMd-aDdBd@dmf/aob5a.d,d*d-b4b7eSc;axb+b.bbcZb0cbfJasdHa/aed+e0cGb/d,btb-b4aWbudpcgdLc=chchd6areOapc0cNb/a;bje/eGaHb5dedOb.a8aNd8aLdLa=a>aIaOaJapb6a+e5azb+cdcfbhc;aOaFdYd6aHaCa@aIaQd8aHa=a.cIbCbMd\\\"\\\",2):f(\\\"\\\"{cycvcocRapcXbocTa;b;bpbgbYdJaGbRanbQaJagbnbcb>dqc5dpbebnbOa8a0c4aJaTa5a+btb5bxbJaQa,c*cRa5a1bzc6aedMa0c3bldjd;aeded8ard5a"));
$write("%s",("6a5aedxb/btbvb2bxb,c1b4b3bxb1b0cocPa8aNapcMagdUc3b|b+b/b2b4arcFbnc4a=a?axbtc4aSbJcPbKckcic+bZb3b-bzcXbqcFb5aMa/ancvc+b+b|byb4a9cVbNa5aRb7cFbnbFbMapb2c.aMaFb.a4a5aJaOa-a-b|b-aeb5aicybHa<b/akc>a>aXb6aOb/a8a6a/apb4a1b.b3bvb4b1b3b2b-b.bvb4anb/aJaPa5a8a4a6apbEb5a5aBb,b9a4apbpbnb8anb4aGa=a:bJacb!\\\"\\\",2):f(\\\"\\\"})23(f\\\"\\\",2):f(\\\"\\\"{#~[2xha=s,y=z,13&X3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'yay,]99999[gnirtS wen=][c n3aea\\\"\\\",2):f(\\\"\\\"{)v]y3b&a(niam diov citats cilbup\\\"\\\",2):f(\\\"\\\"{RQ ssalcz4rfa cdlnl3c/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avajm4bdateg@3doa2 kcats timil.v3dga]; V);"));
$write("%s",("Q4aC3ecaL[b5aX4hha dohtem?3e;4nga repus&3ecaRQ@3cgassalc.<5joa(=:s;0=:c=:i;)|4ajaerudecorp/3fqa(tnirp.biL.oken\\\"\\\",2):f(\\\"\\\"{.3bianoitcnufR6\\\"\\\",2):f(\\\"\\\"{sa(rtStup=niam^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",22):f(\\\"\\\"\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"\\\"\\\",35):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2):f(\\\"\\\"{#v3mja51(f\\\"\\\",2):f(\\\"\\\"{#,4353(ga13(f\\\"\\\",2):f(\\\"\\\"{#j4[j4boa(etirw.z;)tuo.N8aba(67b~auptuOPIZG.piz.litu.avaj wen=zG4Zka30341(f\\\"\\\",2):f(\\\"\\\"{#tm4[m4c5aR0Z0Z/512152353/2/2166263=4/3141726??:1518191:1/@4[@4cda"));
$write("%s",("*6 Q5[p4dea1312^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'5[w8[$5ofa41310r4[r4c7=[B>[j4[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6pma(amirpmi oicy4[(5[j4hma++]371[]591[?6[?6cpani;RQ omtirogla\\\"\\\",2):f(\\\"\\\"{4[\\\"\\\",2):f(\\\"\\\"{4cCa;t:\\\"\\\",2):f(\\\"\\\"}%%%%\\\"\\\",2):f(\\\"\\\"}fi\\\"\\\",2):f(\\\"\\\"}*-84\\\"\\\",2):f(\\\"\\\"})48361(f\\\"\\\",2):f(\\\"\\\"{#]i[\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}+17\\\"\\\",2):f(\\\"\\\"{<84.;i:-i602\\\"\\\",2):f(\\\"\\\""));
$write("%s",("{;i:911\\\"\\\",2):f(\\\"\\\"{;j:632*7[ra116(f\\\"\\\",2):f(\\\"\\\"{#(tnirP.tmfIIcfacnuf;&4[&4bdatmfn4[n4cgaropmi;ILagagakcap~4Zea5102T6dbapD6[r4cba-l4[l4bpatnirp tesn\\\"\\\",2):f(\\\"\\\"})420aEaka etalpmet.r8[ma99(f\\\"\\\",2):f(\\\"\\\"{#(ntnire8[ia974(f\\\"\\\",2):f(\\\"\\\"{#fp4[ga^64^\\\"\\\",2):f(\\\"\\\"})32u9awa,s(llAetirW;)(resUtxeTOPada=:s%8[ba9#8eo4[ia9(f\\\"\\\",2):f(\\\"\\\"{#S Cm4[-Eaca&(y5[ga9(f\\\"\\\",2):f(\\\"\\\"{# .6[.6[.6oiaRQ margo&5[t4cjaS D : ; R-5[6L[j4[j4o%6[k4aqa. EPYT B C : ; Az4[56[j4[j4nka)*,*(ETIRW/6[J7chaA B : ;s4[s4aba [2cr4[*5dia: ^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' ohce3B[EYaeastupLRcdatniy4/ca0"));
$write("%s",("153.ea%%%%m4[m4[53ipaparwyyon noitpoz4023[230ca(nRO.%a7(f\\\"\\\",2):f(\\\"\\\"{#(etirwf:oin\\\"\\\",2):f(\\\"\\\"})4(f\\\"\\\",2):f(\\\"\\\"{#>-)_(niamp3cvP)ka(f\\\"\\\",2):f(\\\"\\\"{# cnirp,L)k;eja.OI[p]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[(3rba@2Wa6;alaM dohtem06x*3c|5aU;cpadiov;oidts.dts 6Yab4kkaenil-etirwb5dva(,^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\""));
$write("%s",(",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'s%^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'(gol.elosnoc;)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'73g\\\"\\\",2):f(\\\"\\\"}a^129^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^"));
$write("%s",("7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' nioj.)1+n(yarrA>-)n(=fI3cwa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"}54,1\\\"\\\",2):f(\\\"\\\"{.^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"# qes-er()|3cH3bba^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"p3lg3fw3hla1% ecalper.j4dea^128^jAc/arts(# pam(]YALPSID^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\""));
$write("%s",("\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NOISIVID ERUDECORPA3cma.RQ .DI-MARGv3g53d|bNOITACIFITNEDI^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"[tac-yzal(s[qesod(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))System.Console.Write($^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Put caffeine \\\"\\\",2):f(\\\"\\\"{(int)c\\\"\\\",2):f(\\\"\\\"} into the mixing bowl.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");M3pva^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Liquify contents ofE3oeaPour^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\"));
$write("%s",("\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3w^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'4e\\\"\\\",2):f(\\\"\\\"{abaking dish.^64^n^64^nServes 164cma\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}/****/e3a^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"),s[999999],*q=s;int main()\\\"\\\",2):f(\\\"\\\"{int n,m;for(;*p;)\\\"\\\",2):f(\\\"\\\"{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>399"));
$write("%s",("9)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\"\\\",2):f(\\\"\\\"}puts(s);return 0;\\\"\\\",2):f(\\\"\\\"}^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(m=1;m<256;m*=2)s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,4,:^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+(c/m%2>0?^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f"));
$write("%s",("(\\\"\\\"\\\\\\\"\\\":^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";f(s);s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4,:,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";\\\"\\\",2):f(\\\"\\\"}f(s+s);for(c:Base64.getDecoder().decode(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"kaAREREX/I0ALn3n5ef6l/Pz8+fnz58/BOf5/7/hEX/OZzM5mCX/OczmZzBPn5+X/OczMznBL/nM5mZzBPu++fP"));
$write("%s",("POc5zngnnOZzOZgnBMGAW7A==^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{c=c<0?256+c:c;for(i=0;i++<3;c/=8)f(c%8);f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8*+8*+,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"@^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");^1^\\\"\\\",4):f(\\\"\\\"'|sed -e^1^\\\"\\\",4):f(\\\"\\\"'s/^16^/^32^/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"/^16^q/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\"));
$write("%s",("\"'s/.*/print ^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^8^nquit/^1^\\\"\\\",4):f(\\\"\\\"'^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",2):f(\\\"\\\"}^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",4):f(\\\"\\\"');\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\").split(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",64):f(\\\"\\\"^\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=1;i<a.length;a[0]+=a[i+1],i+=2)\\\"\\\",2):f(\\\"\\\"{a[0]+=\\\"\\\",25):f(\\\"\\\"\\"));
$write("%s",("\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",89):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".repeat(Integer.parseInt(a[i]));\\\"\\\",2):f(\\\"\\\"}System.out.print(a[0]);\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"J\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+a)OD\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"while(!=(S:length)0)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans c(S:read)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\"));
$write("%s",("\"\\\"\\\\\\\"\\\"D(c:to-integer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 35 39\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 24 149\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"interp:library\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"afnix-sio\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans o(afnix:sio:OutputTerm)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"o:write B\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");end;\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",1):f(\\\"\\\"nsys.exit 0'}\\\\\\\"\\\")\\\"\\\",0)]]></xsl:template></xsl:stylesheet>\\\":s.WriteByte(Asc(c)):Next:End Sub:End Module\")\nput=s\nprint\nqa!"));
end endmodule